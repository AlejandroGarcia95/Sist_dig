library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.includes.all;

-- Componente hardcodeado para inicializar la memoria
-- lógica del Cordic con 510 puntitos x,y,z que representan
-- un tetraedro.

entity init_hardcoded_3d is
   generic (COORD_N: natural := 16; ADDR_N: natural := 12; CANT_PUNTOS : natural := 510);
   port(
      x_out: out std_logic_vector(COORD_N-1 downto 0);
	  y_out: out std_logic_vector(COORD_N-1 downto 0);
	  z_out: out std_logic_vector(COORD_N-1 downto 0);  
	  addr_x: out std_logic_vector(ADDR_N-1 downto 0);
	  addr_y: out std_logic_vector(ADDR_N-1 downto 0);
	  addr_z: out std_logic_vector(ADDR_N-1 downto 0);
	  done: out std_logic;
	  cant_ptos: out std_logic_vector(ADDR_N-1 downto 0);
	  clk: in std_logic
   );
end init_hardcoded_3d;

architecture init_hardcoded_3d_arq of init_hardcoded_3d is
	signal cont_ena: std_logic := '1';
	signal termine: std_logic := '0';
	signal cuenta: std_logic_vector(ADDR_N-1 downto 0);
	type COORDENADAS is array (CANT_PUNTOS-1 downto 0) of std_logic_vector(COORD_N-1 downto 0);	
						                       

--	signal valores_y: COORDENADAS := ("0000000000000000", "0000000001000000", "0000000010000000", "0000000011000001", "0000000100000001", "0000000101000001", "0000000110000010", "0000000111000010", "0000001000000010", "0000001001000011", "0000001010000011", "0000001011000100", "0000001100000100", "0000001101000100", "0000001110000101", "0000001111000101", "0000010000000101", "0000010001000110", "0000010010000110", "0000010011000110", "0000010100000111", "0000010101000111", "0000010110001000", "0000010111001000", "0000011000001000", "0000011001001001", "0000011010001001", "0000011011001001", "0000011100001010", "0000011101001010", "0000011110001010", "0000011111001011", "0000100000001011", "0000100001001100", "0000100010001100", "0000100011001100", "0000100100001101", "0000100101001101", "0000100110001101", "0000100111001110", "0000101000001110", "0000101001001110", "0000101010001111", "0000101011001111", "0000101100010000", "0000101101010000", "0000101110010000", "0000101111010001", "0000110000010001", "0000110001010001", "0000110010010010", "0000110011010010", "0000110100010011", "0000110101010011", "0000110110010011", "0000110111010100", "0000111000010100", "0000111001010100", "0000111010010101", "0000111011010101", "0000111100010101", "0000111101010110", "0000111110010110", "0000111111010111", "0001000000010111", "0001000001010111", "0001000010011000", "0001000011011000", "0001000100011000", "0001000101011001", "0001000110011001", "0001000111011001", "0001001000011010", "0001001001011010", "0001001010011011", "0001001011011011", "0001001100011011", "0001001101011100", "0001001110011100", "0001001111011100", "0001010000011101", "0001010001011101", "0001010010011101", "0001010011011110", "0001010100011110", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000010101", "0000000000101010", "0000000001000000", "0000000001010101", "0000000001101011", "0000000010000000", "0000000010010110", "0000000010101011", "0000000011000001", "0000000011010110", "0000000011101100", "0000000100000001", "0000000100010110", "0000000100101100", "0000000101000001", "0000000101010111", "0000000101101100", "0000000110000010", "0000000110010111", "0000000110101101", "0000000111000010", "0000000111011000", "0000000111101101", "0000001000000010", "0000001000011000", "0000001000101101", "0000001001000011", "0000001001011000", "0000001001101110", "0000001010000011", "0000001010011001", "0000001010101110", "0000001011000100", "0000001011011001", "0000001011101110", "0000001100000100", "0000001100011001", "0000001100101111", "0000001101000100", "0000001101011010", "0000001101101111", "0000001110000101", "0000001110011010", "0000001110110000", "0000001111000101", "0000001111011010", "0000001111110000", "0000010000000101", "0000010000011011", "0000010000110000", "0000010001000110", "0000010001011011", "0000010001110001", "0000010010000110", "0000010010011100", "0000010010110001", "0000010011000110", "0000010011011100", "0000010011110001", "0000010100000111", "0000010100011100", "0000010100110010", "0000010101000111", "0000010101011101", "0000010101110010", "0000010110001000", "0000010110011101", "0000010110110010", "0000010111001000", "0000010111011101", "0000010111110011", "0000011000001000", "0000011000011110", "0000011000110011", "0000011001001001", "0000011001011110", "0000011001110100", "0000011010001001", "0000011010011110", "0000011010110100", "0000011011001001", "0000011011011111", "0000011011110100", "0000011100001010", "0001010100011110", "0001010011011110", "0001010010011101", "0001010001011101", "0001010000011101", "0001001111011100", "0001001110011100", "0001001101011100", "0001001100011011", "0001001011011011", "0001001010011011", "0001001001011010", "0001001000011010", "0001000111011001", "0001000110011001", "0001000101011001", "0001000100011000", "0001000011011000", "0001000010011000", "0001000001010111", "0001000000010111", "0000111111010111", "0000111110010110", "0000111101010110", "0000111100010101", "0000111011010101", "0000111010010101", "0000111001010100", "0000111000010100", "0000110111010100", "0000110110010011", "0000110101010011", "0000110100010011", "0000110011010010", "0000110010010010", "0000110001010001", "0000110000010001", "0000101111010001", "0000101110010000", "0000101101010000", "0000101100010000", "0000101011001111", "0000101010001111", "0000101001001110", "0000101000001110", "0000100111001110", "0000100110001101", "0000100101001101", "0000100100001101", "0000100011001100", "0000100010001100", "0000100001001100", "0000100000001011", "0000011111001011", "0000011110001010", "0000011101001010", "0000011100001010", "0000011011001001", "0000011010001001", "0000011001001001", "0000011000001000", "0000010111001000", "0000010110001000", "0000010101000111", "0000010100000111", "0000010011000110", "0000010010000110", "0000010001000110", "0000010000000101", "0000001111000101", "0000001110000101", "0000001101000100", "0000001100000100", "0000001011000100", "0000001010000011", "0000001001000011", "0000001000000010", "0000000111000010", "0000000110000010", "0000000101000001", "0000000100000001", "0000000011000001", "0000000010000000", "0000000001000000", "0000000000000000", "0001010100011110", "0001010011110011", "0001010011001000", "0001010010011101", "0001010001110011", "0001010001001000", "0001010000011101", "0001001111110010", "0001001111000111", "0001001110011100", "0001001101110001", "0001001101000110", "0001001100011011", "0001001011110000", "0001001011000101", "0001001010011011", "0001001001110000", "0001001001000101", "0001001000011010", "0001000111101111", "0001000111000100", "0001000110011001", "0001000101101110", "0001000101000011", "0001000100011000", "0001000011101101", "0001000011000011", "0001000010011000", "0001000001101101", "0001000001000010", "0001000000010111", "0000111111101100", "0000111111000001", "0000111110010110", "0000111101101011", "0000111101000000", "0000111100010101", "0000111011101011", "0000111011000000", "0000111010010101", "0000111001101010", "0000111000111111", "0000111000010100", "0000110111101001", "0000110110111110", "0000110110010011", "0000110101101000", "0000110100111101", "0000110100010011", "0000110011101000", "0000110010111101", "0000110010010010", "0000110001100111", "0000110000111100", "0000110000010001", "0000101111100110", "0000101110111011", "0000101110010000", "0000101101100101", "0000101100111011", "0000101100010000", "0000101011100101", "0000101010111010", "0000101010001111", "0000101001100100", "0000101000111001", "0000101000001110", "0000100111100011", "0000100110111000", "0000100110001101", "0000100101100010", "0000100100111000", "0000100100001101", "0000100011100010", "0000100010110111", "0000100010001100", "0000100001100001", "0000100000110110", "0000100000001011", "0000011111100000", "0000011110110101", "0000011110001010", "0000011101100000", "0000011100110101", "0000011100001010", "0000000000000000", "0000000000010101", "0000000000101010", "0000000001000000", "0000000001010101", "0000000001101011", "0000000010000000", "0000000010010110", "0000000010101011", "0000000011000001", "0000000011010110", "0000000011101100", "0000000100000001", "0000000100010110", "0000000100101100", "0000000101000001", "0000000101010111", "0000000101101100", "0000000110000010", "0000000110010111", "0000000110101101", "0000000111000010", "0000000111011000", "0000000111101101", "0000001000000010", "0000001000011000", "0000001000101101", "0000001001000011", "0000001001011000", "0000001001101110", "0000001010000011", "0000001010011001", "0000001010101110", "0000001011000100", "0000001011011001", "0000001011101110", "0000001100000100", "0000001100011001", "0000001100101111", "0000001101000100", "0000001101011010", "0000001101101111", "0000001110000101", "0000001110011010", "0000001110110000", "0000001111000101", "0000001111011010", "0000001111110000", "0000010000000101", "0000010000011011", "0000010000110000", "0000010001000110", "0000010001011011", "0000010001110001", "0000010010000110", "0000010010011100", "0000010010110001", "0000010011000110", "0000010011011100", "0000010011110001", "0000010100000111", "0000010100011100", "0000010100110010", "0000010101000111", "0000010101011101", "0000010101110010", "0000010110001000", "0000010110011101", "0000010110110010", "0000010111001000", "0000010111011101", "0000010111110011", "0000011000001000", "0000011000011110", "0000011000110011", "0000011001001001", "0000011001011110", "0000011001110100", "0000011010001001", "0000011010011110", "0000011010110100", "0000011011001001", "0000011011011111", "0000011011110100", "0000011100001010");
--	signal valores_z: COORDENADAS := ("0000000000000000", "0000000000100101", "0000000001001010", "0000000001101111", "0000000010010100", "0000000010111001", "0000000011011110", "0000000100000011", "0000000100101000", "0000000101001101", "0000000101110010", "0000000110010111", "0000000110111100", "0000000111100001", "0000001000000110", "0000001000101011", "0000001001010000", "0000001001110110", "0000001010011011", "0000001011000000", "0000001011100101", "0000001100001010", "0000001100101111", "0000001101010100", "0000001101111001", "0000001110011110", "0000001111000011", "0000001111101000", "0000010000001101", "0000010000110010", "0000010001010111", "0000010001111100", "0000010010100001", "0000010011000110", "0000010011101100", "0000010100010001", "0000010100110110", "0000010101011011", "0000010110000000", "0000010110100101", "0000010111001010", "0000010111101111", "0000011000010100", "0000011000111001", "0000011001011110", "0000011010000011", "0000011010101000", "0000011011001101", "0000011011110010", "0000011100010111", "0000011100111100", "0000011101100010", "0000011110000111", "0000011110101100", "0000011111010001", "0000011111110110", "0000100000011011", "0000100001000000", "0000100001100101", "0000100010001010", "0000100010101111", "0000100011010100", "0000100011111001", "0000100100011110", "0000100101000011", "0000100101101000", "0000100110001101", "0000100110110010", "0000100111011000", "0000100111111101", "0000101000100010", "0000101001000111", "0000101001101100", "0000101010010001", "0000101010110110", "0000101011011011", "0000101100000000", "0000101100100101", "0000101101001010", "0000101101101111", "0000101110010100", "0000101110111001", "0000101111011110", "0000110000000011", "0000110000101000", "0000000000000000", "0000000001001010", "0000000010010100", "0000000011011110", "0000000100101000", "0000000101110010", "0000000110111100", "0000001000000110", "0000001001010000", "0000001010011011", "0000001011100101", "0000001100101111", "0000001101111001", "0000001111000011", "0000010000001101", "0000010001010111", "0000010010100001", "0000010011101100", "0000010100110110", "0000010110000000", "0000010111001010", "0000011000010100", "0000011001011110", "0000011010101000", "0000011011110010", "0000011100111100", "0000011110000111", "0000011111010001", "0000100000011011", "0000100001100101", "0000100010101111", "0000100011111001", "0000100101000011", "0000100110001101", "0000100111011000", "0000101000100010", "0000101001101100", "0000101010110110", "0000101100000000", "0000101101001010", "0000101110010100", "0000101111011110", "0000110000101000", "0000110001110011", "0000110010111101", "0000110100000111", "0000110101010001", "0000110110011011", "0000110111100101", "0000111000101111", "0000111001111001", "0000111011000100", "0000111100001110", "0000111101011000", "0000111110100010", "0000111111101100", "0001000000110110", "0001000010000000", "0001000011001010", "0001000100010100", "0001000101011111", "0001000110101001", "0001000111110011", "0001001000111101", "0001001010000111", "0001001011010001", "0001001100011011", "0001001101100101", "0001001110110000", "0001001111111010", "0001010001000100", "0001010010001110", "0001010011011000", "0001010100100010", "0001010101101100", "0001010110110110", "0001011000000000", "0001011001001011", "0001011010010101", "0001011011011111", "0001011100101001", "0001011101110011", "0001011110111101", "0001100000000111", "0001100001010001", "0000000000000000", "0000000000100101", "0000000001001010", "0000000001101111", "0000000010010100", "0000000010111001", "0000000011011110", "0000000100000011", "0000000100101000", "0000000101001101", "0000000101110010", "0000000110010111", "0000000110111100", "0000000111100001", "0000001000000110", "0000001000101011", "0000001001010000", "0000001001110110", "0000001010011011", "0000001011000000", "0000001011100101", "0000001100001010", "0000001100101111", "0000001101010100", "0000001101111001", "0000001110011110", "0000001111000011", "0000001111101000", "0000010000001101", "0000010000110010", "0000010001010111", "0000010001111100", "0000010010100001", "0000010011000110", "0000010011101100", "0000010100010001", "0000010100110110", "0000010101011011", "0000010110000000", "0000010110100101", "0000010111001010", "0000010111101111", "0000011000010100", "0000011000111001", "0000011001011110", "0000011010000011", "0000011010101000", "0000011011001101", "0000011011110010", "0000011100010111", "0000011100111100", "0000011101100010", "0000011110000111", "0000011110101100", "0000011111010001", "0000011111110110", "0000100000011011", "0000100001000000", "0000100001100101", "0000100010001010", "0000100010101111", "0000100011010100", "0000100011111001", "0000100100011110", "0000100101000011", "0000100101101000", "0000100110001101", "0000100110110010", "0000100111011000", "0000100111111101", "0000101000100010", "0000101001000111", "0000101001101100", "0000101010010001", "0000101010110110", "0000101011011011", "0000101100000000", "0000101100100101", "0000101101001010", "0000101101101111", "0000101110010100", "0000101110111001", "0000101111011110", "0000110000000011", "0000110000101000", "0000110000101000", "0000110001001110", "0000110001110011", "0000110010011000", "0000110010111101", "0000110011100010", "0000110100000111", "0000110100101100", "0000110101010001", "0000110101110110", "0000110110011011", "0000110111000000", "0000110111100101", "0000111000001010", "0000111000101111", "0000111001010100", "0000111001111001", "0000111010011110", "0000111011000100", "0000111011101001", "0000111100001110", "0000111100110011", "0000111101011000", "0000111101111101", "0000111110100010", "0000111111000111", "0000111111101100", "0001000000010001", "0001000000110110", "0001000001011011", "0001000010000000", "0001000010100101", "0001000011001010", "0001000011101111", "0001000100010100", "0001000100111010", "0001000101011111", "0001000110000100", "0001000110101001", "0001000111001110", "0001000111110011", "0001001000011000", "0001001000111101", "0001001001100010", "0001001010000111", "0001001010101100", "0001001011010001", "0001001011110110", "0001001100011011", "0001001101000000", "0001001101100101", "0001001110001010", "0001001110110000", "0001001111010101", "0001001111111010", "0001010000011111", "0001010001000100", "0001010001101001", "0001010010001110", "0001010010110011", "0001010011011000", "0001010011111101", "0001010100100010", "0001010101000111", "0001010101101100", "0001010110010001", "0001010110110110", "0001010111011011", "0001011000000000", "0001011000100110", "0001011001001011", "0001011001110000", "0001011010010101", "0001011010111010", "0001011011011111", "0001011100000100", "0001011100101001", "0001011101001110", "0001011101110011", "0001011110011000", "0001011110111101", "0001011111100010", "0001100000000111", "0001100000101100", "0001100001010001", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0000110000101000", "0001100001010001", "0001100000101100", "0001100000000111", "0001011111100010", "0001011110111101", "0001011110011000", "0001011101110011", "0001011101001110", "0001011100101001", "0001011100000100", "0001011011011111", "0001011010111010", "0001011010010101", "0001011001110000", "0001011001001011", "0001011000100110", "0001011000000000", "0001010111011011", "0001010110110110", "0001010110010001", "0001010101101100", "0001010101000111", "0001010100100010", "0001010011111101", "0001010011011000", "0001010010110011", "0001010010001110", "0001010001101001", "0001010001000100", "0001010000011111", "0001001111111010", "0001001111010101", "0001001110110000", "0001001110001010", "0001001101100101", "0001001101000000", "0001001100011011", "0001001011110110", "0001001011010001", "0001001010101100", "0001001010000111", "0001001001100010", "0001001000111101", "0001001000011000", "0001000111110011", "0001000111001110", "0001000110101001", "0001000110000100", "0001000101011111", "0001000100111010", "0001000100010100", "0001000011101111", "0001000011001010", "0001000010100101", "0001000010000000", "0001000001011011", "0001000000110110", "0001000000010001", "0000111111101100", "0000111111000111", "0000111110100010", "0000111101111101", "0000111101011000", "0000111100110011", "0000111100001110", "0000111011101001", "0000111011000100", "0000111010011110", "0000111001111001", "0000111001010100", "0000111000101111", "0000111000001010", "0000110111100101", "0000110111000000", "0000110110011011", "0000110101110110", "0000110101010001", "0000110100101100", "0000110100000111", "0000110011100010", "0000110010111101", "0000110010011000", "0000110001110011", "0000110001001110", "0000110000101000");
--	signal valores_x: COORDENADAS := ("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000111100", "0000000001111000", "0000000010110101", "0000000011110001", "0000000100101110", "0000000101101010", "0000000110100111", "0000000111100011", "0000001000100000", "0000001001011100", "0000001010011001", "0000001011010101", "0000001100010010", "0000001101001110", "0000001110001010", "0000001111000111", "0000010000000011", "0000010001000000", "0000010001111100", "0000010010111001", "0000010011110101", "0000010100110010", "0000010101101110", "0000010110101011", "0000010111100111", "0000011000100100", "0000011001100000", "0000011010011101", "0000011011011001", "0000011100010101", "0000011101010010", "0000011110001110", "0000011111001011", "0000100000000111", "0000100001000100", "0000100010000000", "0000100010111101", "0000100011111001", "0000100100110110", "0000100101110010", "0000100110101111", "0000100111101011", "0000101000100111", "0000101001100100", "0000101010100000", "0000101011011101", "0000101100011001", "0000101101010110", "0000101110010010", "0000101111001111", "0000110000001011", "0000110001001000", "0000110010000100", "0000110011000001", "0000110011111101", "0000110100111010", "0000110101110110", "0000110110110010", "0000110111101111", "0000111000101011", "0000111001101000", "0000111010100100", "0000111011100001", "0000111100011101", "0000111101011010", "0000111110010110", "0000111111010011", "0001000000001111", "0001000001001100", "0001000010001000", "0001000011000100", "0001000100000001", "0001000100111101", "0001000101111010", "0001000110110110", "0001000111110011", "0001001000101111", "0001001001101100", "0001001010101000", "0001001011100101", "0001001100100001", "0001001101011110", "0001001110011010", "0001001111010111", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000111100", "0000000001111000", "0000000010110101", "0000000011110001", "0000000100101110", "0000000101101010", "0000000110100111", "0000000111100011", "0000001000100000", "0000001001011100", "0000001010011001", "0000001011010101", "0000001100010010", "0000001101001110", "0000001110001010", "0000001111000111", "0000010000000011", "0000010001000000", "0000010001111100", "0000010010111001", "0000010011110101", "0000010100110010", "0000010101101110", "0000010110101011", "0000010111100111", "0000011000100100", "0000011001100000", "0000011010011101", "0000011011011001", "0000011100010101", "0000011101010010", "0000011110001110", "0000011111001011", "0000100000000111", "0000100001000100", "0000100010000000", "0000100010111101", "0000100011111001", "0000100100110110", "0000100101110010", "0000100110101111", "0000100111101011", "0000101000100111", "0000101001100100", "0000101010100000", "0000101011011101", "0000101100011001", "0000101101010110", "0000101110010010", "0000101111001111", "0000110000001011", "0000110001001000", "0000110010000100", "0000110011000001", "0000110011111101", "0000110100111010", "0000110101110110", "0000110110110010", "0000110111101111", "0000111000101011", "0000111001101000", "0000111010100100", "0000111011100001", "0000111100011101", "0000111101011010", "0000111110010110", "0000111111010011", "0001000000001111", "0001000001001100", "0001000010001000", "0001000011000100", "0001000100000001", "0001000100111101", "0001000101111010", "0001000110110110", "0001000111110011", "0001001000101111", "0001001001101100", "0001001010101000", "0001001011100101", "0001001100100001", "0001001101011110", "0001001110011010", "0001001111010111", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000");											   
	signal valores_x: COORDENADAS := ("0000000000000000", "0001000000000000", "0000000000000000", "0001000000000000", "0000000000000000", "0001000000000000", "0000000000000000", "0001000000000000", "0000000000000000");
	signal valores_y: COORDENADAS := ("0000000000000000", "0000000000000000", "0001000000000000", "0001000000000000", "0000000000000000", "0000000000000000", "0001000000000000", "0001000000000000", "0000000000000000");
	signal valores_z: COORDENADAS := ("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000","0001000000000000", "0001000000000000", "0001000000000000", "0001000000000000", "0000000000000000");
begin													                       
	process(clk)
	begin
		if rising_edge(clk) then
			x_out <= valores_x(to_integer(unsigned(cuenta)));
			y_out <= valores_y(to_integer(unsigned(cuenta)));
			z_out <= valores_z(to_integer(unsigned(cuenta)));
			addr_x <= cuenta;
			addr_y <= cuenta;
			addr_z <= cuenta; -- Ojo aquí !! Strong assumption!
		end if;
 		if (to_integer(unsigned(cuenta)) = CANT_PUNTOS-1) then 
 			cont_ena <= '0';
 			termine <= '1';
 		else
 			cont_ena <= '1';
 			termine <= '0';
 		end if;
	end process;

	myCounter: contador
		generic map(N => ADDR_N)
		port map (clk, '0', cont_ena, cuenta);

	flipflop: ffd
		port map(clk, '0', '1', termine, done);
		
	cant_ptos <= std_logic_vector(to_unsigned(CANT_PUNTOS, ADDR_N));

end init_hardcoded_3d_arq;