library IEEE;
use IEEE.std_logic_1164.all;
use work.includes_TP2.all;

entity video_log_tb is
end;

architecture beh of video_log_tb is

begin

end beh;