library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Char_ROM is
    generic(
        N: integer:= 6;
        M: integer:= 3;
        W: integer:= 8
    );
    port(
        char_address: in std_logic_vector(5 downto 0);
        font_row, font_col: in std_logic_vector(M-1 downto 0);
        rom_out: out std_logic
    );
end;

architecture p of Char_ROM is
    subtype tipoLinea is std_logic_vector(0 to W-1);

    type char is array(0 to W-1) of tipoLinea;
     
    constant NUM_0: char:= (
                                "00111100",
                                "01100110",
                                "01101110",
                                "01111110",
                                "01110110",
                                "01100110",
                                "00111100",
                                "00000000"
                        );  
						
    constant NUM_1: char:= (
                                "00000000",
                                "00001000",
                                "00011000",
                                "00101000",
                                "00001000",
                                "00001000",
                                "00011100",
                                "00000000"
                        );
					     
    constant NUM_2: char:= (
                                "00000000",
                                "00111100",
                                "00110110",
                                "00000110",
                                "00001100",
                                "00011000",
                                "00111110",
                                "00000000"
                        );  
						
    constant NUM_3: char:= (
                                "00000000",
                                "00111100",
                                "00000110",
                                "00011110",
                                "00000110",
                                "00000110",
                                "00111100",
                                "00000000"
                        );
     
    constant NUM_4: char:= (
                                "00001000",
                                "00011000",
                                "00101000",
                                "01001000",
                                "01111100",
                                "00001000",
                                "00001000",
                                "00000000"
                        );  
						
    constant NUM_5: char:= (
                                "00000000",
                                "00111100",
                                "00100000",
                                "00110000",
                                "00001100",
                                "00001100",
                                "00111000",
                                "00000000"
                        );
					     
    constant NUM_6: char:= (
                                "00000000",
                                "00111100",
                                "01100000",
                                "01111100",
                                "01100110",
                                "01100110",
                                "00111100",
                                "00000000"
                        );  
						
    constant NUM_7: char:= (
                                "00000000",
                                "00111110",
                                "00100110",
                                "00001100",
                                "00001000",
                                "00011000",
                                "00011000",
                                "00000000"
                        );     
    constant NUM_8: char:= (
                                "00111100",
                                "01100110",
                                "01100110",
                                "01111110",
                                "01100110",
                                "01100110",
                                "00111100",
                                "00000000"
                        );  
						
    constant NUM_9: char:= (
                                "00000000",
                                "00111100",
                                "01100110",
                                "01100110",								
                                "00111110",								
                                "00000110",
                                "00111100",
                                "00000000"
                        );
					     
    constant V: char:= (
                                "00000000",
                                "01000010",
                                "01100110",
                                "01100110",
                                "01100110",
                                "00111100",
                                "00011000",
                                "00000000"
                        );  
						
    constant COMMA: char:= (
                                "00000000",
                                "00000000",
		                        "00000000",
                                "00000000",
                                "00000000",
                                "00001000",
		                        "00011000",
                                "00010000"
                        );
	
					
	constant A: char:= (
                                "00011000",
                                "00111100",
                                "01100110",
                                "01100110",
                                "01111110",
                                "01100110",
                                "01100110",
                                "00000000"
                        );
    constant B: char:= (
                                "01111100",
                                "01100110",
                                "01100110",
                                "01111100",
                                "01100110",
                                "01100110",
                                "01111100",
                                "00000000"
                        );
    constant C: char:= (
                                "00111110",
                                "01100011",
                                "01100000",
                                "01100000",
                                "01100000",
                                "01100011",
                                "00111110",
                                "00000000"
                        );

    constant D: char:= (
                                "01111100",
                                "01100110",
                                "01100011",
                                "01100011",
                                "01100011",
                                "01100110",
                                "01111100",
                                "00000000"
                        );

    constant E: char:= (
                                "01111110",
                                "01100000",
                                "01100000",
                                "01111000",
                                "01100000",
                                "01100000",
                                "01111110",
                                "00000000"
                        );

    constant F: char:= (
                                "01111110",
                                "01100000",
                                "01100000",
                                "01111000",
                                "01100000",
                                "01100000",
                                "01100000",
                                "00000000"
                        );

    constant G: char:= (
                                "00111100",
                                "01100010",
                                "01100000",
                                "01101110",
                                "01100110",
                                "01100110",
                                "00111100",
                                "00000000"
                        );

    constant H: char:= (
                                "01100110",
                                "01100110",
                                "01100110",
                                "01111110",
                                "01100110",
                                "01100110",
                                "01100110",
                                "00000000"
                        );
                        
    constant N_Char: char:= (
                             "01100110",
                             "01100110",
                             "01110110",
                             "01110110",
                             "01101110",
                             "01101110",
                             "01100110",
                             "00000000"
                     );
                        
    constant O: char:= (
                                "00111100",
                                "01100110",
                                "01100110",
                                "01100110",
                                "01100110",
                                "01100110",
                                "00111100",
                                "00000000"
                        );
                        
    constant Err: char:= (
                                "00000000",
                                "01111110",
                                "01111110",
                                "01100110",
                                "01100110",
                                "01111110",
                                "01111110",
                                "00000000"
                        );
                        

    type memo is array(0 to 255) of tipoLinea;
    signal RAM: memo:= (
                                0 => NUM_0(0), 1 => NUM_0(1), 2 => NUM_0(2), 3 => NUM_0(3), 4 => NUM_0(4), 5 => NUM_0(5), 6 => NUM_0(6), 7 => NUM_0(7),
                                8 => NUM_1(0), 9 => NUM_1(1), 10 => NUM_1(2), 11 => NUM_1(3), 12 => NUM_1(4), 13 => NUM_1(5), 14 => NUM_1(6), 15 => NUM_1(7),
                                16 => NUM_2(0), 17 => NUM_2(1), 18 => NUM_2(2), 19 => NUM_2(3), 20 => NUM_2(4), 21 => NUM_2(5), 22 => NUM_2(6), 23 => NUM_2(7),
                                24 => NUM_3(0), 25 => NUM_3(1), 26 => NUM_3(2), 27 => NUM_3(3), 28 => NUM_3(4), 29 => NUM_3(5), 30 => NUM_3(6), 31 => NUM_3(7),
                                32 => NUM_4(0), 33 => NUM_4(1), 34 => NUM_4(2), 35 => NUM_4(3), 36 => NUM_4(4), 37 => NUM_4(5), 38 => NUM_4(6), 39 => NUM_4(7),
                                40 => NUM_5(0), 41 => NUM_5(1), 42 => NUM_5(2), 43 => NUM_5(3), 44 => NUM_5(4), 45 => NUM_5(5), 46 => NUM_5(6), 47 => NUM_5(7),
                                48 => NUM_6(0), 49 => NUM_6(1), 50 => NUM_6(2), 51 => NUM_6(3), 52 => NUM_6(4), 53 => NUM_6(5), 54 => NUM_6(6), 55 => NUM_6(7),
                                56 => NUM_7(0), 57 => NUM_7(1), 58 => NUM_7(2), 59 => NUM_7(3), 60 => NUM_7(4), 61 => NUM_7(5), 62 => NUM_7(6), 63 => NUM_7(7),
                                64 => NUM_8(0), 65 => NUM_8(1), 66 => NUM_8(2), 67 => NUM_8(3), 68 => NUM_8(4), 69 => NUM_8(5), 70 => NUM_8(6), 71 => NUM_8(7),
                                72 => NUM_9(0), 73 => NUM_9(1), 74 => NUM_9(2), 75 => NUM_9(3), 76 => NUM_9(4), 77 => NUM_9(5), 78 => NUM_9(6), 79 => NUM_9(7),
								80 => V(0), 81 => V(1), 82 => V(2), 83 => V(3), 84 => V(4), 85 => V(5), 86 => V(6), 87 => V(7),
								88 => COMMA(0), 89 => COMMA(1), 90=> COMMA(2), 91 => COMMA(3), 92 => COMMA(4), 93 => COMMA(5), 94 => COMMA(6), 95 => COMMA(7),
                           
                                96 => Err(0), 97 => Err(1), 98 => Err(2), 99 => Err(3), 100 => Err(4), 101 => Err(5), 102 => Err(6), 103 => Err(7),
                                104 to 255 => "00000000"
                            );

    signal char_addr_aux: std_logic_vector(8 downto 0);
    
begin

    char_addr_aux <= char_address & font_row;
    rom_out <= RAM(conv_integer(char_addr_aux))(conv_integer(font_col));

end;
